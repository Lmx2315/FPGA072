module versiya_fpga072 (
	output [47:0] data	
);

reg [47:0] ver_data=48'h290320211706;//29-03-2021 17-06

endmodule